* /media/camilo/data/workspaces/personal_projects/the_wah_pedal/pcb_kicad/wah_pedal.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Wed 16 Aug 2017 06:24:05 PM JST

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
R1  /Input Net-_C1-Pad2_ 68kR		
C1  Net-_C1-Pad1_ Net-_C1-Pad2_ 0.01uF		
R2  Net-_C4-Pad2_ Net-_C1-Pad1_ 1.5kR		
R4  Net-_R4-Pad1_ Net-_Q1-Pade_ 470R		
R3  Net-_C3-Pad2_ Net-_R3-Pad2_ 22kR		
L1  Net-_C4-Pad2_ Net-_C2-Pad1_ 500mH		
R5  Net-_C2-Pad1_ Net-_C3-Pad2_ 470kR		
R6  Net-_C4-Pad2_ Net-_C2-Pad1_ 33kR		
R7  Net-_C2-Pad2_ Net-_C2-Pad1_ 82kR		
C4  Net-_C4-Pad1_ Net-_C4-Pad2_ 0.01uF		
R9  Net-_C3-Pad2_ Net-_C5-Pad1_ 470kR		
C5  Net-_C5-Pad1_ Net-_C5-Pad2_ 0.22uF		
C3  /Output Net-_C3-Pad2_ 0.22uF		
R10  Net-_Q2-Padc_ Net-_R10-Pad2_ 1kR		
R11  Net-_R11-Pad1_ Net-_C4-Pad1_ 10kR		
R8  Net-_R8-Pad1_ /Output Net-_C5-Pad2_ 100kR		
Q1  Net-_C1-Pad1_ Net-_C3-Pad2_ Net-_Q1-Pade_ Q-NPN-BEC		
Q2  Net-_C5-Pad1_ Net-_Q2-Padc_ Net-_C4-Pad1_ Q-NPN-BEC		
C2  Net-_C2-Pad1_ Net-_C2-Pad2_ 4.7uF		
P1  /Input 01X01		
P2  /Output CONN_01X01		
P4  Net-_P4-Pad1_ 01X01		
P3  Net-_P3-Pad1_ 01X01		

.end
